library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mixColumnTB is
end entity;

architecture tb_arch of mixColumnTB is
    -- Constants
    constant CLOCK_PERIOD : time := 10 ns;
    
    -- Signals
    signal clk : std_logic := '0';
    signal i_block : std_logic_vector(127 downto 0) := (others => '0');
    signal valid_i : std_logic := '0';
    signal valid_o : std_logic;
    signal o_block : std_logic_vector(127 downto 0);

    -- Component instantiation
    component mixColumn
        port (
            clk     : in std_logic;
            i_block : in std_logic_vector(127 downto 0);
            o_block : out std_logic_vector(127 downto 0);
            valid_i : in std_logic;
            valid_o : out std_logic
        );
    end component;

begin
    -- DUT (Device Under Test) instantiation
    DUT: mixColumn
    port map (
        clk => clk,
        i_block => i_block,
        o_block => o_block,
        valid_i => valid_i,
        valid_o => valid_o
    );

    -- Clock process
    clk_process: process
    begin
        while now < 1000 ns loop
            clk <= '0';
            wait for CLOCK_PERIOD / 2;
            clk <= '1';
            wait for CLOCK_PERIOD / 2;
        end loop;
        wait;
    end process;

    -- Stimulus process
    stimulus: process
    begin
        -- Wait for initializations

        -- Input data
        i_block <= x"25252525252525252525252525252525"; -- Example input data
         wait for 10 ns;
        valid_i <= '1'; -- Set valid input

        wait for 100 ns; -- Wait for some time

        -- Additional stimuli can be added here as needed

        wait;
    end process;

end tb_arch;
