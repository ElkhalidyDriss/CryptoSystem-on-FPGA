-- ==========================================================================
-- Project        : AES-128
-- File           : multiplier2x2.vhd
-- Authors        : Meziani EL-Houcine 
--                  Elkhalidy Driss
--
-- Date           : May 2024
-- Version        : 1.0
-- 
-- Description    : Implementation of the a multiplier in GF(2^2) to be used in the shiftRows calculations.
-- 
-- ==========================================================================


library ieee;
use ieee.std_logic_1164.all;

--Entity for a 2x2 multiplier in GF(2^2)
entity mutliplier2x2 is
port (  i_data1 : in std_logic_vector(1 downto 0);   --input data 1 in GF(2^2)
        i_data2 : in std_logic_vector(1 downto 0);   --input data 2 in GF(2^2)
        o_data : out std_logic_vector(1 downto 0));  --output data result in GF(2^2) of multiplication of the two inputs
end entity;


architecture mutliplier2x2Arch of mutliplier2x2 is

begin
o_data(1) <= (i_data1(0) and i_data2(1)) xor (i_data1(1) and (i_data2(0) xor i_data2(1)));
o_data(0) <= (i_data1(1) and i_data2(1)) xor (i_data2(0) and i_data1(0));
end architecture;