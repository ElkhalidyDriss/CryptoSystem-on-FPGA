library ieee;
use ieee.std_logic_1164.all;


entity subByte is 
port(
     i_data : in std_logic_vector(7 downto 0); --input data in GF(2^8)
     o_data : out std_logic_vector(7 downto 0)-- output data
);
end entity;

architecture subByteArch of subByte is 
begin
process(i_data)
begin
case i_data is
          when x"00" => o_data <= x"63";
          when x"01" => o_data <= x"7c";
          when x"02" => o_data <= x"77";
          when x"03" => o_data <= x"7b";
          when x"04" => o_data <= x"f2";
          when x"05" => o_data <= x"6b";
          when x"06" => o_data <= x"6f";
          when x"07" => o_data <= x"c5";
          when x"08" => o_data <= x"30";
          when x"09" => o_data <= x"01";
          when x"0a" => o_data <= x"67";
          when x"0b" => o_data <= x"2b";
          when x"0c" => o_data <= x"fe";
          when x"0d" => o_data <= x"d7";
          when x"0e" => o_data <= x"ab";
          when x"0f" => o_data <= x"76";
          when x"10" => o_data <= x"ca";
          when x"11" => o_data <= x"82";
          when x"12" => o_data <= x"c9";
          when x"13" => o_data <= x"7d";
          when x"14" => o_data <= x"fa";
          when x"15" => o_data <= x"59";
          when x"16" => o_data <= x"47";
          when x"17" => o_data <= x"f0";
          when x"18" => o_data <= x"ad";
          when x"19" => o_data <= x"d4";
          when x"1a" => o_data <= x"a2";
          when x"1b" => o_data <= x"af";
          when x"1c" => o_data <= x"9c";
          when x"1d" => o_data <= x"a4";
          when x"1e" => o_data <= x"72";
          when x"1f" => o_data <= x"c0";
          when x"20" => o_data <= x"b7";
          when x"21" => o_data <= x"fd";
          when x"22" => o_data <= x"93";
          when x"23" => o_data <= x"26";
          when x"24" => o_data <= x"36";
          when x"25" => o_data <= x"3f";
          when x"26" => o_data <= x"f7";
          when x"27" => o_data <= x"cc";
          when x"28" => o_data <= x"34";
          when x"29" => o_data <= x"a5";
          when x"2a" => o_data <= x"e5";
          when x"2b" => o_data <= x"f1";
          when x"2c" => o_data <= x"71";
          when x"2d" => o_data <= x"d8";
          when x"2e" => o_data <= x"31";
          when x"2f" => o_data <= x"15";
          when x"30" => o_data <= x"04";
          when x"31" => o_data <= x"c7";
          when x"32" => o_data <= x"23";
          when x"33" => o_data <= x"c3";
          when x"34" => o_data <= x"18";
          when x"35" => o_data <= x"96";
          when x"36" => o_data <= x"05";
          when x"37" => o_data <= x"9a";
          when x"38" => o_data <= x"07";
          when x"39" => o_data <= x"12";
          when x"3a" => o_data <= x"80";
          when x"3b" => o_data <= x"e2";
          when x"3c" => o_data <= x"eb";
          when x"3d" => o_data <= x"27";
          when x"3e" => o_data <= x"b2";
          when x"3f" => o_data <= x"75";
          when x"40" => o_data <= x"09";
          when x"41" => o_data <= x"83";
          when x"42" => o_data <= x"2c";
          when x"43" => o_data <= x"1a";
          when x"44" => o_data <= x"1b";
          when x"45" => o_data <= x"6e";
          when x"46" => o_data <= x"5a";
          when x"47" => o_data <= x"a0";
          when x"48" => o_data <= x"52";
          when x"49" => o_data <= x"3b";
          when x"4a" => o_data <= x"d6";
          when x"4b" => o_data <= x"b3";
          when x"4c" => o_data <= x"29";
          when x"4d" => o_data <= x"e3";
          when x"4e" => o_data <= x"2f";
          when x"4f" => o_data <= x"84";
          when x"50" => o_data <= x"53";
          when x"51" => o_data <= x"d1";
          when x"52" => o_data <= x"00";
          when x"53" => o_data <= x"ed";
          when x"54" => o_data <= x"20";
          when x"55" => o_data <= x"fc";
          when x"56" => o_data <= x"b1";
          when x"57" => o_data <= x"5b";
          when x"58" => o_data <= x"6a";
          when x"59" => o_data <= x"cb";
          when x"5a" => o_data <= x"be";
          when x"5b" => o_data <= x"39";
          when x"5c" => o_data <= x"4a";
          when x"5d" => o_data <= x"4c";
          when x"5e" => o_data <= x"58";
          when x"5f" => o_data <= x"cf";
          when x"60" => o_data <= x"d0";
          when x"61" => o_data <= x"ef";
          when x"62" => o_data <= x"aa";
          when x"63" => o_data <= x"fb";
          when x"64" => o_data <= x"43";
          when x"65" => o_data <= x"4d";
          when x"66" => o_data <= x"33";
          when x"67" => o_data <= x"85";
          when x"68" => o_data <= x"45";
          when x"69" => o_data <= x"f9";
          when x"6a" => o_data <= x"02";
          when x"6b" => o_data <= x"7f";
          when x"6c" => o_data <= x"50";
          when x"6d" => o_data <= x"3c";
          when x"6e" => o_data <= x"9f";
          when x"6f" => o_data <= x"a8";
          when x"70" => o_data <= x"51";
          when x"71" => o_data <= x"a3";
          when x"72" => o_data <= x"40";
          when x"73" => o_data <= x"8f";
          when x"74" => o_data <= x"92";
          when x"75" => o_data <= x"9d";
          when x"76" => o_data <= x"38";
          when x"77" => o_data <= x"f5";
          when x"78" => o_data <= x"bc";
          when x"79" => o_data <= x"b6";
          when x"7a" => o_data <= x"da";
          when x"7b" => o_data <= x"21";
          when x"7c" => o_data <= x"10";
          when x"7d" => o_data <= x"ff";
          when x"7e" => o_data <= x"f3";
          when x"7f" => o_data <= x"d2";
          when x"80" => o_data <= x"cd";
          when x"81" => o_data <= x"0c";
          when x"82" => o_data <= x"13";
          when x"83" => o_data <= x"ec";
          when x"84" => o_data <= x"5f";
          when x"85" => o_data <= x"97";
          when x"86" => o_data <= x"44";
          when x"87" => o_data <= x"17";
          when x"88" => o_data <= x"c4";
          when x"89" => o_data <= x"a7";
          when x"8a" => o_data <= x"7e";
          when x"8b" => o_data <= x"3d";
          when x"8c" => o_data <= x"64";
          when x"8d" => o_data <= x"5d";
          when x"8e" => o_data <= x"19";
          when x"8f" => o_data <= x"73";
          when x"90" => o_data <= x"60";
          when x"91" => o_data <= x"81";
          when x"92" => o_data <= x"4f";
          when x"93" => o_data <= x"dc";
          when x"94" => o_data <= x"22";
          when x"95" => o_data <= x"2a";
          when x"96" => o_data <= x"90";
          when x"97" => o_data <= x"88";
          when x"98" => o_data <= x"46";
          when x"99" => o_data <= x"ee";
          when x"9a" => o_data <= x"b8";
          when x"9b" => o_data <= x"14";
          when x"9c" => o_data <= x"de";
          when x"9d" => o_data <= x"5e";
          when x"9e" => o_data <= x"0b";
          when x"9f" => o_data <= x"db";
          when x"a0" => o_data <= x"e0";
          when x"a1" => o_data <= x"32";
          when x"a2" => o_data <= x"3a";
          when x"a3" => o_data <= x"0a";
          when x"a4" => o_data <= x"49";
          when x"a5" => o_data <= x"06";
          when x"a6" => o_data <= x"24";
          when x"a7" => o_data <= x"5c";
          when x"a8" => o_data <= x"c2";
          when x"a9" => o_data <= x"d3";
          when x"aa" => o_data <= x"ac";
          when x"ab" => o_data <= x"62";
          when x"ac" => o_data <= x"91";
          when x"ad" => o_data <= x"95";
          when x"ae" => o_data <= x"e4";
          when x"af" => o_data <= x"79";
          when x"b0" => o_data <= x"e7";
          when x"b1" => o_data <= x"c8";
          when x"b2" => o_data <= x"37";
          when x"b3" => o_data <= x"6d";
          when x"b4" => o_data <= x"8d";
          when x"b5" => o_data <= x"d5";
          when x"b6" => o_data <= x"4e";
          when x"b7" => o_data <= x"a9";
          when x"b8" => o_data <= x"6c";
          when x"b9" => o_data <= x"56";
          when x"ba" => o_data <= x"f4";
          when x"bb" => o_data <= x"ea";
          when x"bc" => o_data <= x"65";
          when x"bd" => o_data <= x"7a";
          when x"be" => o_data <= x"ae";
          when x"bf" => o_data <= x"08";
          when x"c0" => o_data <= x"ba";
          when x"c1" => o_data <= x"78";
          when x"c2" => o_data <= x"25";
          when x"c3" => o_data <= x"2e";
          when x"c4" => o_data <= x"1c";
          when x"c5" => o_data <= x"a6";
          when x"c6" => o_data <= x"b4";
          when x"c7" => o_data <= x"c6";
          when x"c8" => o_data <= x"e8";
          when x"c9" => o_data <= x"dd";
          when x"ca" => o_data <= x"74";
          when x"cb" => o_data <= x"1f";
          when x"cc" => o_data <= x"4b";
          when x"cd" => o_data <= x"bd";
          when x"ce" => o_data <= x"8b";
          when x"cf" => o_data <= x"8a";
          when x"d0" => o_data <= x"70";
          when x"d1" => o_data <= x"3e";
          when x"d2" => o_data <= x"b5";
          when x"d3" => o_data <= x"66";
          when x"d4" => o_data <= x"48";
          when x"d5" => o_data <= x"03";
          when x"d6" => o_data <= x"f6";
          when x"d7" => o_data <= x"0e";
          when x"d8" => o_data <= x"61";
          when x"d9" => o_data <= x"35";
          when x"da" => o_data <= x"57";
          when x"db" => o_data <= x"b9";
          when x"dc" => o_data <= x"86";
          when x"dd" => o_data <= x"c1";
          when x"de" => o_data <= x"1d";
          when x"df" => o_data <= x"9e";
          when x"e0" => o_data <= x"e1";
          when x"e1" => o_data <= x"f8";
          when x"e2" => o_data <= x"98";
          when x"e3" => o_data <= x"11";
          when x"e4" => o_data <= x"69";
          when x"e5" => o_data <= x"d9";
          when x"e6" => o_data <= x"8e";
          when x"e7" => o_data <= x"94";
          when x"e8" => o_data <= x"9b";
          when x"e9" => o_data <= x"1e";
          when x"ea" => o_data <= x"87";
          when x"eb" => o_data <= x"e9";
          when x"ec" => o_data <= x"ce";
          when x"ed" => o_data <= x"55";
          when x"ee" => o_data <= x"28";
          when x"ef" => o_data <= x"df";
          when x"f0" => o_data <= x"8c";
          when x"f1" => o_data <= x"a1";
          when x"f2" => o_data <= x"89";
          when x"f3" => o_data <= x"0d";
          when x"f4" => o_data <= x"bf";
          when x"f5" => o_data <= x"e6";
          when x"f6" => o_data <= x"42";
          when x"f7" => o_data <= x"68";
          when x"f8" => o_data <= x"41";
          when x"f9" => o_data <= x"99";
          when x"fa" => o_data <= x"2d";
          when x"fb" => o_data <= x"0f";
          when x"fc" => o_data <= x"b0";
          when x"fd" => o_data <= x"54";
          when x"fe" => o_data <= x"bb";
          when x"ff" => o_data <= x"16";
 when others => null;
end case;
end process;
end architecture;