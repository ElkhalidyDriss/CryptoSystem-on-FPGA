library ieee;
use ieee.std_logic_1164.all;


entity subByte is 
port(
     i_data : in std_logic_vector(7 downto 0); --input data
     o_data : out std_logic_vector(7 downto 0)-- output data
);
end entity;

architecture subByteArch of subByte is 


begin



end architecture;